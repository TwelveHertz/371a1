module display (register, Hex);
	input [31:0] register;
	output reg [6:0] Hex; 
	

endmodule