module storeOperand (current, store);
	input [11:0] current;
	output [11:0] store;
	
	assign store = current;
		
endmodule